`define ADDR_ACQ_CR                    4'h0
`define ACQ_CR_START_OFFSET 0
`define ACQ_CR_START 32'h00000001
`define ACQ_CR_READY_OFFSET 1
`define ACQ_CR_READY 32'h00000002
`define ADDR_ACQ_ADDR                  4'h4
`define ADDR_ACQ_DATA                  4'h8
