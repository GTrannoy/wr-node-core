`define ADDR_TOF_MINTREV               4'h0
`define ADDR_TOF_MAXTREV               4'h4
`define ADDR_TOF_CTRL                  4'h8
`define TOF_CTRL_WRLTCY_OFFSET 0
`define TOF_CTRL_WRLTCY 32'h000fffff
`define TOF_CTRL_GMARGIN_OFFSET 24
`define TOF_CTRL_GMARGIN 32'h03000000
`define TOF_CTRL_GWIDTH_OFFSET 26
`define TOF_CTRL_GWIDTH 32'h0c000000
