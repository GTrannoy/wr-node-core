`define ADDR_WRN_CPU_CSR_APP_ID        7'h0
`define ADDR_WRN_CPU_CSR_RESET         7'h4
`define ADDR_WRN_CPU_CSR_ENABLE        7'h8
`define ADDR_WRN_CPU_CSR_UADDR         7'hc
`define WRN_CPU_CSR_UADDR_ADDR_OFFSET 0
`define WRN_CPU_CSR_UADDR_ADDR 32'h000fffff
`define ADDR_WRN_CPU_CSR_CORE_SEL      7'h10
`define ADDR_WRN_CPU_CSR_CORE_COUNT    7'h14
`define ADDR_WRN_CPU_CSR_CORE_MEMSIZE  7'h18
`define ADDR_WRN_CPU_CSR_UDATA         7'h1c
`define ADDR_WRN_CPU_CSR_DBG_JTAG      7'h20
`define WRN_CPU_CSR_DBG_JTAG_JDATA_OFFSET 0
`define WRN_CPU_CSR_DBG_JTAG_JDATA 32'h000000ff
`define WRN_CPU_CSR_DBG_JTAG_JADDR_OFFSET 8
`define WRN_CPU_CSR_DBG_JTAG_JADDR 32'h00000700
`define WRN_CPU_CSR_DBG_JTAG_RSTN_OFFSET 16
`define WRN_CPU_CSR_DBG_JTAG_RSTN 32'h00010000
`define WRN_CPU_CSR_DBG_JTAG_TCK_OFFSET 17
`define WRN_CPU_CSR_DBG_JTAG_TCK 32'h00020000
`define WRN_CPU_CSR_DBG_JTAG_UPDATE_OFFSET 18
`define WRN_CPU_CSR_DBG_JTAG_UPDATE 32'h00040000
`define ADDR_WRN_CPU_CSR_DBG_MSG       7'h24
`define WRN_CPU_CSR_DBG_MSG_DATA_OFFSET 0
`define WRN_CPU_CSR_DBG_MSG_DATA 32'h000000ff
`define ADDR_WRN_CPU_CSR_DBG_POLL      7'h28
`define WRN_CPU_CSR_DBG_POLL_READY_OFFSET 0
`define WRN_CPU_CSR_DBG_POLL_READY 32'h000000ff
`define ADDR_WRN_CPU_CSR_DBG_IMSK      7'h2c
`define WRN_CPU_CSR_DBG_IMSK_ENABLE_OFFSET 0
`define WRN_CPU_CSR_DBG_IMSK_ENABLE 32'h000000ff
`define ADDR_WRN_CPU_CSR_SMEM_OP       7'h30
`define ADDR_WRN_CPU_CSR_TPU_CSR       7'h34
`define WRN_CPU_CSR_TPU_CSR_PRESENT_OFFSET 0
`define WRN_CPU_CSR_TPU_CSR_PRESENT 32'h00000001
`define WRN_CPU_CSR_TPU_CSR_ENABLE_OFFSET 1
`define WRN_CPU_CSR_TPU_CSR_ENABLE 32'h00000002
`define WRN_CPU_CSR_TPU_CSR_FORCE_START_OFFSET 2
`define WRN_CPU_CSR_TPU_CSR_FORCE_START 32'h00000004
`define WRN_CPU_CSR_TPU_CSR_READY_OFFSET 3
`define WRN_CPU_CSR_TPU_CSR_READY 32'h00000008
`define WRN_CPU_CSR_TPU_CSR_PROBE_COUNT_OFFSET 4
`define WRN_CPU_CSR_TPU_CSR_PROBE_COUNT 32'h000001f0
`define WRN_CPU_CSR_TPU_CSR_PROBE_SEL_OFFSET 9
`define WRN_CPU_CSR_TPU_CSR_PROBE_SEL 32'h00003e00
`define ADDR_WRN_CPU_CSR_TPU_PROBE_CSR 7'h38
`define WRN_CPU_CSR_TPU_PROBE_CSR_PC_OFFSET 0
`define WRN_CPU_CSR_TPU_PROBE_CSR_PC 32'h00ffffff
`define WRN_CPU_CSR_TPU_PROBE_CSR_CORE_ID_OFFSET 24
`define WRN_CPU_CSR_TPU_PROBE_CSR_CORE_ID 32'h0f000000
`define WRN_CPU_CSR_TPU_PROBE_CSR_ACTION_OFFSET 28
`define WRN_CPU_CSR_TPU_PROBE_CSR_ACTION 32'hf0000000
`define ADDR_WRN_CPU_CSR_TPU_BUF_COUNT 7'h3c
`define ADDR_WRN_CPU_CSR_TPU_BUF_SIZE  7'h40
`define ADDR_WRN_CPU_CSR_TPU_BUF_ADDR  7'h44
`define ADDR_WRN_CPU_CSR_TPU_BUF_DATA  7'h48
`define WRN_CPU_CSR_TPU_BUF_DATA_ID_OFFSET 0
`define WRN_CPU_CSR_TPU_BUF_DATA_ID 32'h0000001f
`define WRN_CPU_CSR_TPU_BUF_DATA_TSTAMP_OFFSET 5
`define WRN_CPU_CSR_TPU_BUF_DATA_TSTAMP 32'hffffffe0
