`define ADDR_D3SS_RSTR                 6'h0
`define D3SS_RSTR_PLL_RST_OFFSET 0
`define D3SS_RSTR_PLL_RST 32'h00000001
`define ADDR_D3SS_TCR                  6'h4
`define D3SS_TCR_WR_LOCK_EN_OFFSET 0
`define D3SS_TCR_WR_LOCK_EN 32'h00000001
`define D3SS_TCR_WR_LOCKED_OFFSET 1
`define D3SS_TCR_WR_LOCKED 32'h00000002
`define D3SS_TCR_WR_TIME_VALID_OFFSET 2
`define D3SS_TCR_WR_TIME_VALID 32'h00000004
`define D3SS_TCR_WR_LINK_OFFSET 3
`define D3SS_TCR_WR_LINK 32'h00000008
`define ADDR_D3SS_GPIOR                6'h8
`define D3SS_GPIOR_PLL_SYS_CS_N_OFFSET 0
`define D3SS_GPIOR_PLL_SYS_CS_N 32'h00000001
`define D3SS_GPIOR_PLL_SYS_RESET_N_OFFSET 1
`define D3SS_GPIOR_PLL_SYS_RESET_N 32'h00000002
`define D3SS_GPIOR_PLL_SCLK_OFFSET 2
`define D3SS_GPIOR_PLL_SCLK 32'h00000004
`define D3SS_GPIOR_PLL_SDIO_OFFSET 3
`define D3SS_GPIOR_PLL_SDIO 32'h00000008
`define D3SS_GPIOR_PLL_SDIO_DIR_OFFSET 4
`define D3SS_GPIOR_PLL_SDIO_DIR 32'h00000010
`define D3SS_GPIOR_PLL_VCXO_RESET_N_OFFSET 5
`define D3SS_GPIOR_PLL_VCXO_RESET_N 32'h00000020
`define D3SS_GPIOR_PLL_VCXO_CS_N_OFFSET 6
`define D3SS_GPIOR_PLL_VCXO_CS_N 32'h00000040
`define D3SS_GPIOR_PLL_VCXO_SDO_OFFSET 7
`define D3SS_GPIOR_PLL_VCXO_SDO 32'h00000080
`define D3SS_GPIOR_ADF_CE_OFFSET 8
`define D3SS_GPIOR_ADF_CE 32'h00000100
`define D3SS_GPIOR_ADF_CLK_OFFSET 9
`define D3SS_GPIOR_ADF_CLK 32'h00000200
`define D3SS_GPIOR_ADF_LE_OFFSET 10
`define D3SS_GPIOR_ADF_LE 32'h00000400
`define D3SS_GPIOR_ADF_DATA_OFFSET 11
`define D3SS_GPIOR_ADF_DATA 32'h00000800
`define D3SS_GPIOR_SERDES_PLL_LOCKED_OFFSET 12
`define D3SS_GPIOR_SERDES_PLL_LOCKED 32'h00001000
`define ADDR_D3SS_CR                   6'hc
`define D3SS_CR_ENABLE_OFFSET 0
`define D3SS_CR_ENABLE 32'h00000001
`define ADDR_D3SS_REC_DELAY_COARSE     6'h10
`define ADDR_D3SS_FREV_TS_SEC          6'h14
`define ADDR_D3SS_FREV_TS_NS           6'h18
`define ADDR_D3SS_FREV_CR              6'h1c
`define D3SS_FREV_CR_VALID_OFFSET 0
`define D3SS_FREV_CR_VALID 32'h00000001
`define D3SS_FREV_CR_READY_OFFSET 1
`define D3SS_FREV_CR_READY 32'h00000002
`define ADDR_D3SS_PHFIFO_R0            6'h20
`define D3SS_PHFIFO_R0_PAYLOAD_OFFSET 0
`define D3SS_PHFIFO_R0_PAYLOAD 32'hffffffff
`define ADDR_D3SS_PHFIFO_CSR           6'h24
`define D3SS_PHFIFO_CSR_FULL_OFFSET 16
`define D3SS_PHFIFO_CSR_FULL 32'h00010000
`define D3SS_PHFIFO_CSR_EMPTY_OFFSET 17
`define D3SS_PHFIFO_CSR_EMPTY 32'h00020000
`define D3SS_PHFIFO_CSR_CLEAR_BUS_OFFSET 18
`define D3SS_PHFIFO_CSR_CLEAR_BUS 32'h00040000
`define D3SS_PHFIFO_CSR_USEDW_OFFSET 0
`define D3SS_PHFIFO_CSR_USEDW 32'h000003ff
