`define ADDR_D3S_TCR                   6'h0
`define D3S_TCR_WR_LOCK_EN_OFFSET 0
`define D3S_TCR_WR_LOCK_EN 32'h00000001
`define D3S_TCR_WR_LOCKED_OFFSET 1
`define D3S_TCR_WR_LOCKED 32'h00000002
`define D3S_TCR_WR TIME VALID_OFFSET 2
`define D3S_TCR_WR TIME VALID 32'h00000004
`define D3S_TCR_WR_LINK_OFFSET 3
`define D3S_TCR_WR_LINK 32'h00000008
`define ADDR_D3S_GPIOR                 6'h4
`define D3S_GPIOR_SI57X_SCL_OFFSET 0
`define D3S_GPIOR_SI57X_SCL 32'h00000001
`define D3S_GPIOR_SI57X_SDA_OFFSET 1
`define D3S_GPIOR_SI57X_SDA 32'h00000002
`define D3S_GPIOR_SPI_CS_ADC_OFFSET 2
`define D3S_GPIOR_SPI_CS_ADC 32'h00000004
`define D3S_GPIOR_SPI_SCK_OFFSET 3
`define D3S_GPIOR_SPI_SCK 32'h00000008
`define D3S_GPIOR_SPI_MOSI_OFFSET 4
`define D3S_GPIOR_SPI_MOSI 32'h00000010
`define D3S_GPIOR_SPI_MISO_OFFSET 5
`define D3S_GPIOR_SPI_MISO 32'h00000020
`define ADDR_D3S_SSR                   6'h8
`define ADDR_D3S_CR                    6'hc
`define D3S_CR_ENABLE_OFFSET 0
`define D3S_CR_ENABLE 32'h00000001
`define ADDR_D3S_RL_ERR_MIN            6'h10
`define ADDR_D3S_RL_ERR_MAX            6'h14
`define ADDR_D3S_RL_LENGTH_MAX         6'h18
`define ADDR_D3S_ADC_R0                6'h1c
`define D3S_ADC_R0_TSTAMP_OFFSET 0
`define D3S_ADC_R0_TSTAMP 32'h0fffffff
`define D3S_ADC_R0_IS_RL_OFFSET 28
`define D3S_ADC_R0_IS_RL 32'h10000000
`define ADDR_D3S_ADC_R1                6'h20
`define D3S_ADC_R1_RL_LENGTH_OFFSET 0
`define D3S_ADC_R1_RL_LENGTH 32'h0000ffff
`define ADDR_D3S_ADC_R2                6'h24
`define D3S_ADC_R2_RL_PHASE_OFFSET 0
`define D3S_ADC_R2_RL_PHASE 32'hffffffff
`define ADDR_D3S_ADC_CSR               6'h28
`define D3S_ADC_CSR_FULL_OFFSET 16
`define D3S_ADC_CSR_FULL 32'h00010000
`define D3S_ADC_CSR_EMPTY_OFFSET 17
`define D3S_ADC_CSR_EMPTY 32'h00020000
`define D3S_ADC_CSR_CLEAR_BUS_OFFSET 18
`define D3S_ADC_CSR_CLEAR_BUS 32'h00040000
`define D3S_ADC_CSR_USEDW_OFFSET 0
`define D3S_ADC_CSR_USEDW 32'h000003ff
