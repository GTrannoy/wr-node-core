`define ADDR_TREVGEN_RM_NEXT_TICK      5'h0
`define ADDR_TREVGEN_LC_NEXT_TICK      5'h4
`define ADDR_TREVGEN_RM_TREV           5'h8
`define ADDR_TREVGEN_LC_TREV           5'hc
`define ADDR_TREVGEN_STROBE_P          5'h10
