`define ADDR_TREVGEN_RM_NEXT_TICK      4'h0
`define ADDR_TREVGEN_RM_TREV           4'h4
`define ADDR_TREVGEN_STROBE_P          4'h8
`define ADDR_TREVGEN_DUMMY             4'hc
`define TREVGEN_DUMMY_DUMMY_OFFSET 0
`define TREVGEN_DUMMY_DUMMY 32'h00000001
