`define ADDR_TDCSERDES_STATUS          4'h0
`define TDCSERDES_STATUS_NOEMPTY_OFFSET 0
`define TDCSERDES_STATUS_NOEMPTY 32'h00000001
`define TDCSERDES_STATUS_OF_OFFSET 1
`define TDCSERDES_STATUS_OF 32'h00000002
`define ADDR_TDCSERDES_CTRL            4'h4
`define TDCSERDES_CTRL_CLR_OFFSET 0
`define TDCSERDES_CTRL_CLR 32'h00000001
`define TDCSERDES_CTRL_CLR_OF_OFFSET 1
`define TDCSERDES_CTRL_CLR_OF 32'h00000002
`define TDCSERDES_CTRL_NEXT_OFFSET 2
`define TDCSERDES_CTRL_NEXT 32'h00000004
`define TDCSERDES_CTRL_FILTER_OFFSET 3
`define TDCSERDES_CTRL_FILTER 32'h00000018
`define ADDR_TDCSERDES_TDC_DATA        4'h8
`define TDCSERDES_TDC_DATA_TDC_DATA_OFFSET 0
`define TDCSERDES_TDC_DATA_TDC_DATA 32'hffffffff
