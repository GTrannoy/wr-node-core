`define ADDR_STDC_STATUS               4'h0
`define STDC_STATUS_EMPTY_OFFSET 0
`define STDC_STATUS_EMPTY 32'h00000001
`define STDC_STATUS_OVF_OFFSET 1
`define STDC_STATUS_OVF 32'h00000002
`define ADDR_STDC_CTRL                 4'h4
`define STDC_CTRL_CLR_OFFSET 0
`define STDC_CTRL_CLR 32'h00000001
`define STDC_CTRL_CLR_OVF_OFFSET 1
`define STDC_CTRL_CLR_OVF 32'h00000002
`define STDC_CTRL_NEXT_OFFSET 2
`define STDC_CTRL_NEXT 32'h00000004
`define STDC_CTRL_FILTER_OFFSET 3
`define STDC_CTRL_FILTER 32'h00000018
`define ADDR_STDC_TDC_DATA             4'h8
